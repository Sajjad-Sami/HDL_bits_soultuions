Exams/m2014 q4i
module top_module (
    output out);
assign out = 1'b0;
endmodule
