//Exams/m2014 q4h
module top_module (
    input in,
    output out);
assign out = in;
endmodule
